library IEEE;
use IEEE.STD_LOGIC_1164.all;

package UMDRISC_PKG is
	CONSTANT INSTR_MEM_WIDTH: INTEGER := 12;
end UMDRISC_PKG;

package body UMDRISC_PKG is

end UMDRISC_PKG;
